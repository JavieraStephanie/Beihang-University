`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:53:43 12/05/2019 
// Design Name: 
// Module Name:    stop 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module stop(
	 input [31:0] ir_d,
	 input [31:0] ir_e,
	 input [31:0] ir_m,
	 output delay
    );


endmodule
